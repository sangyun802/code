module Datapath(

);
    reg [15:0] pc, read_data1, read_data2, ALUout, memorydata;

endmodule